`timescale 1ns / 1ps


module audio(
    input clock

    );
    
    always @(posedge clock)
    begin
    
    
    
    end
endmodule
